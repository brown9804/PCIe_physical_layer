// Belinda Brown Ramírez
// Mayo, 2020
// timna.brown@ucr.ac.cr

// 						&


/////////////////////////////////////////////////////////////////////////////////
// Company: U.C.R EIE
// Engineer: Brandon Esquivel Molina
//
//////////////////////////////////////////////////////////////////////////////////

`timescale 	1ns				/ 1ps
`include "./lib/cmos_cells.v"
`include "./src/demux1x2_behav.v"
`include "./syn/demux1x2_behav_syn.v"
`include "./testers/t_demux12.v"



module TestBench;


/// 						COLOCAR EL REAL

endmodule
